CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
12
10 555 Timer~
219 877 312 0 8 17
0 18 19 20 21 22 23 24 25
0
0 0 4944 0
3 555
-11 -36 10 -28
2 U5
-7 -46 7 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 512 1 0 0 0
1 U
5130 0 0
2
43529.9 0
0
7 Ground~
168 1145 61 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
43529.9 1
0
2 +V
167 294 256 0 1 3
0 7
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.89883e-315 0
0
7 Pulser~
4 96 305 0 10 12
0 26 27 8 28 0 0 5 5 3
8
0
0 0 6704 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3421 0 0
2
5.89883e-315 5.26354e-315
0
9 CC 7-Seg~
183 1146 149 0 17 19
10 15 14 13 12 11 10 9 29 2
1 1 1 0 0 0 0 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8157 0 0
2
5.89883e-315 5.30499e-315
0
9 2-In AND~
219 703 211 0 3 22
0 16 4 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5572 0 0
2
5.89883e-315 5.32571e-315
0
9 2-In AND~
219 523 200 0 3 22
0 6 5 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8901 0 0
2
5.89883e-315 5.34643e-315
0
6 74112~
219 781 335 0 7 32
0 7 17 8 17 7 30 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
7361 0 0
2
5.89883e-315 5.3568e-315
0
6 74112~
219 617 333 0 7 32
0 7 16 8 16 7 4 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
4747 0 0
2
5.89883e-315 5.36716e-315
0
6 74112~
219 441 336 0 7 32
0 7 6 8 6 7 31 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
972 0 0
2
5.89883e-315 5.37752e-315
0
6 74112~
219 294 336 0 7 32
0 7 7 8 7 7 32 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3472 0 0
2
5.89883e-315 5.38788e-315
0
6 74LS48
188 1015 282 0 14 29
0 3 4 5 6 33 34 9 10 11
12 13 14 15 35
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.89883e-315 5.39306e-315
0
38
0 0 3 0 0 4096 0 0 0 4 0 2
827 299
851 299
6 0 4 0 0 12288 0 9 0 0 5 4
647 315
641 315
641 315
671 315
1 9 2 0 0 12416 0 2 5 0 0 4
1145 69
1145 84
1146 84
1146 107
7 1 3 0 0 16512 0 8 12 0 0 6
805 299
828 299
828 357
938 357
938 246
983 246
0 2 4 0 0 8336 0 0 12 30 0 5
671 297
671 367
947 367
947 255
983 255
0 3 5 0 0 8320 0 0 12 28 0 5
483 300
483 380
957 380
957 264
983 264
0 4 6 0 0 8320 0 0 12 38 0 5
333 300
333 391
966 391
966 273
983 273
0 1 7 0 0 8192 0 0 3 25 0 4
256 300
256 273
294 273
294 265
1 0 7 0 0 0 0 3 0 0 13 2
294 265
294 265
0 0 7 0 0 4096 0 0 0 13 16 2
355 265
355 356
1 1 7 0 0 8192 0 9 8 0 0 4
617 270
617 265
781 265
781 272
1 1 7 0 0 8320 0 10 9 0 0 4
441 273
441 265
617 265
617 270
1 1 7 0 0 0 0 11 10 0 0 4
294 273
294 265
441 265
441 273
5 5 7 0 0 0 0 9 8 0 0 4
617 345
617 356
781 356
781 347
5 5 7 0 0 0 0 10 9 0 0 4
441 348
441 356
617 356
617 345
5 5 7 0 0 0 0 11 10 0 0 4
294 348
294 356
441 356
441 348
3 0 8 0 0 8192 0 4 0 0 35 4
120 296
140 296
140 410
242 410
7 7 9 0 0 4224 0 12 5 0 0 3
1047 246
1161 246
1161 185
8 6 10 0 0 4224 0 12 5 0 0 3
1047 255
1155 255
1155 185
9 5 11 0 0 4224 0 12 5 0 0 3
1047 264
1149 264
1149 185
10 4 12 0 0 4224 0 12 5 0 0 3
1047 273
1143 273
1143 185
11 3 13 0 0 8320 0 12 5 0 0 3
1047 282
1137 282
1137 185
12 2 14 0 0 8320 0 12 5 0 0 3
1047 291
1131 291
1131 185
13 1 15 0 0 8320 0 12 5 0 0 3
1047 300
1125 300
1125 185
4 2 7 0 0 0 0 11 11 0 0 4
270 318
256 318
256 300
270 300
2 0 16 0 0 4096 0 9 0 0 27 2
593 297
548 297
0 4 16 0 0 4224 0 0 9 29 0 3
548 200
548 315
593 315
2 7 5 0 0 0 0 7 10 0 0 4
499 209
492 209
492 300
465 300
3 1 16 0 0 12416 0 7 6 0 0 4
544 200
548 200
548 202
679 202
2 7 4 0 0 0 0 6 9 0 0 3
679 220
679 297
641 297
2 0 17 0 0 4096 0 8 0 0 32 2
757 299
733 299
3 4 17 0 0 8320 0 6 8 0 0 4
724 211
733 211
733 317
757 317
3 0 8 0 0 0 0 9 0 0 35 3
587 306
554 306
554 410
3 0 8 0 0 0 0 10 0 0 35 3
411 309
397 309
397 410
3 3 8 0 0 12416 0 11 8 0 0 6
264 309
242 309
242 410
702 410
702 308
751 308
1 0 6 0 0 0 0 7 0 0 37 3
499 191
367 191
367 300
4 0 6 0 0 0 0 10 0 0 38 3
417 318
367 318
367 300
7 2 6 0 0 0 0 11 10 0 0 2
318 300
417 300
3
-27 0 0 0 700 0 0 0 0 3 2 1 34
16 Arial Unicode MS
0 0 0 35
282 84 931 137
300 93 912 130
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
-27 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
318 9 497 56
332 18 482 49
10 BS CpE 1-B
-27 0 0 0 700 255 0 0 0 3 2 1 18
10 Constantia
0 0 0 17
5 7 273 54
23 16 254 49
17 Jumamoy, Davee S.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
